// ============================================================
// Exponential Lookup Table (for Softmax)
// Input  : 16-bit signed (Q8.7) in range [-8, 0]
// Output : 12-bit unsigned Q1.11 (e^x)
// ============================================================

module exp_lut (
    input  logic signed [15:0] input_q8_7,    // Q8.7 signed input
    output logic [11:0] output_q1_11   // Q1.11 unsigned output
);

    logic [7:0] lut_index;  // 8-bit index for 256-entry LUT
    // Convert Q8.7 input to LUT index
    always_comb begin
        // Q8.7 range [-8, 0] maps to indices [0, 255]
        // -8.0 in Q8.7 = 16'hFC00 = -1024
        // 0.0 in Q8.7  = 16'h0000 = 0

        if (input_q8_7 >= 16'shFC00 && input_q8_7 < 16'sh0000) begin
            // Map [-1024, 0] to [0, 255]
            // index = (input + 1024) / 4
            lut_index = (input_q8_7 + 16'sh0400) >>> 2;  // Add 1024, then divide by 4
        end else if (input_q8_7 < 16'shFC00) begin
            lut_index = 8'h00;  // Clamp to minimum (most negative)
        end else begin
            lut_index = 8'hFF;  // Clamp to maximum (zero)
        end
    end
	

    always_comb begin
        case (lut_index)
            8'h00: output_q1_11 = 12'h000; // e^(-8.000) = 0.000335
            8'h01: output_q1_11 = 12'h000; // e^(-7.969) = 0.000346
            8'h02: output_q1_11 = 12'h000; // e^(-7.937) = 0.000357
            8'h03: output_q1_11 = 12'h000; // e^(-7.906) = 0.000369
            8'h04: output_q1_11 = 12'h000; // e^(-7.875) = 0.000380
            8'h05: output_q1_11 = 12'h000; // e^(-7.843) = 0.000392
            8'h06: output_q1_11 = 12'h000; // e^(-7.812) = 0.000405
            8'h07: output_q1_11 = 12'h000; // e^(-7.780) = 0.000418
            8'h08: output_q1_11 = 12'h000; // e^(-7.749) = 0.000431
            8'h09: output_q1_11 = 12'h000; // e^(-7.718) = 0.000445
            8'h0A: output_q1_11 = 12'h000; // e^(-7.686) = 0.000459
            8'h0B: output_q1_11 = 12'h000; // e^(-7.655) = 0.000474
            8'h0C: output_q1_11 = 12'h001; // e^(-7.624) = 0.000489
            8'h0D: output_q1_11 = 12'h001; // e^(-7.592) = 0.000504
            8'h0E: output_q1_11 = 12'h001; // e^(-7.561) = 0.000520
            8'h0F: output_q1_11 = 12'h001; // e^(-7.529) = 0.000537
            8'h10: output_q1_11 = 12'h001; // e^(-7.498) = 0.000554
            8'h11: output_q1_11 = 12'h001; // e^(-7.467) = 0.000572
            8'h12: output_q1_11 = 12'h001; // e^(-7.435) = 0.000590
            8'h13: output_q1_11 = 12'h001; // e^(-7.404) = 0.000609
            8'h14: output_q1_11 = 12'h001; // e^(-7.373) = 0.000628
            8'h15: output_q1_11 = 12'h001; // e^(-7.341) = 0.000648
            8'h16: output_q1_11 = 12'h001; // e^(-7.310) = 0.000669
            8'h17: output_q1_11 = 12'h001; // e^(-7.278) = 0.000690
            8'h18: output_q1_11 = 12'h001; // e^(-7.247) = 0.000712
            8'h19: output_q1_11 = 12'h001; // e^(-7.216) = 0.000735
            8'h1A: output_q1_11 = 12'h001; // e^(-7.184) = 0.000758
            8'h1B: output_q1_11 = 12'h001; // e^(-7.153) = 0.000783
            8'h1C: output_q1_11 = 12'h001; // e^(-7.122) = 0.000807
            8'h1D: output_q1_11 = 12'h001; // e^(-7.090) = 0.000833
            8'h1E: output_q1_11 = 12'h001; // e^(-7.059) = 0.000860
            8'h1F: output_q1_11 = 12'h001; // e^(-7.027) = 0.000887
            8'h20: output_q1_11 = 12'h001; // e^(-6.996) = 0.000915
            8'h21: output_q1_11 = 12'h001; // e^(-6.965) = 0.000945
            8'h22: output_q1_11 = 12'h001; // e^(-6.933) = 0.000975
            8'h23: output_q1_11 = 12'h002; // e^(-6.902) = 0.001006
            8'h24: output_q1_11 = 12'h002; // e^(-6.871) = 0.001038
            8'h25: output_q1_11 = 12'h002; // e^(-6.839) = 0.001071
            8'h26: output_q1_11 = 12'h002; // e^(-6.808) = 0.001105
            8'h27: output_q1_11 = 12'h002; // e^(-6.776) = 0.001140
            8'h28: output_q1_11 = 12'h002; // e^(-6.745) = 0.001177
            8'h29: output_q1_11 = 12'h002; // e^(-6.714) = 0.001214
            8'h2A: output_q1_11 = 12'h002; // e^(-6.682) = 0.001253
            8'h2B: output_q1_11 = 12'h002; // e^(-6.651) = 0.001293
            8'h2C: output_q1_11 = 12'h002; // e^(-6.620) = 0.001334
            8'h2D: output_q1_11 = 12'h002; // e^(-6.588) = 0.001376
            8'h2E: output_q1_11 = 12'h002; // e^(-6.557) = 0.001420
            8'h2F: output_q1_11 = 12'h003; // e^(-6.525) = 0.001466
            8'h30: output_q1_11 = 12'h003; // e^(-6.494) = 0.001512
            8'h31: output_q1_11 = 12'h003; // e^(-6.463) = 0.001561
            8'h32: output_q1_11 = 12'h003; // e^(-6.431) = 0.001610
            8'h33: output_q1_11 = 12'h003; // e^(-6.400) = 0.001662
            8'h34: output_q1_11 = 12'h003; // e^(-6.369) = 0.001715
            8'h35: output_q1_11 = 12'h003; // e^(-6.337) = 0.001769
            8'h36: output_q1_11 = 12'h003; // e^(-6.306) = 0.001826
            8'h37: output_q1_11 = 12'h003; // e^(-6.275) = 0.001884
            8'h38: output_q1_11 = 12'h003; // e^(-6.243) = 0.001944
            8'h39: output_q1_11 = 12'h004; // e^(-6.212) = 0.002006
            8'h3A: output_q1_11 = 12'h004; // e^(-6.180) = 0.002070
            8'h3B: output_q1_11 = 12'h004; // e^(-6.149) = 0.002136
            8'h3C: output_q1_11 = 12'h004; // e^(-6.118) = 0.002204
            8'h3D: output_q1_11 = 12'h004; // e^(-6.086) = 0.002274
            8'h3E: output_q1_11 = 12'h004; // e^(-6.055) = 0.002346
            8'h3F: output_q1_11 = 12'h004; // e^(-6.024) = 0.002421
            8'h40: output_q1_11 = 12'h005; // e^(-5.992) = 0.002498
            8'h41: output_q1_11 = 12'h005; // e^(-5.961) = 0.002578
            8'h42: output_q1_11 = 12'h005; // e^(-5.929) = 0.002660
            8'h43: output_q1_11 = 12'h005; // e^(-5.898) = 0.002745
            8'h44: output_q1_11 = 12'h005; // e^(-5.867) = 0.002832
            8'h45: output_q1_11 = 12'h005; // e^(-5.835) = 0.002923
            8'h46: output_q1_11 = 12'h006; // e^(-5.804) = 0.003016
            8'h47: output_q1_11 = 12'h006; // e^(-5.773) = 0.003112
            8'h48: output_q1_11 = 12'h006; // e^(-5.741) = 0.003211
            8'h49: output_q1_11 = 12'h006; // e^(-5.710) = 0.003313
            8'h4A: output_q1_11 = 12'h007; // e^(-5.678) = 0.003419
            8'h4B: output_q1_11 = 12'h007; // e^(-5.647) = 0.003528
            8'h4C: output_q1_11 = 12'h007; // e^(-5.616) = 0.003640
            8'h4D: output_q1_11 = 12'h007; // e^(-5.584) = 0.003756
            8'h4E: output_q1_11 = 12'h007; // e^(-5.553) = 0.003876
            8'h4F: output_q1_11 = 12'h008; // e^(-5.522) = 0.004000
            8'h50: output_q1_11 = 12'h008; // e^(-5.490) = 0.004127
            8'h51: output_q1_11 = 12'h008; // e^(-5.459) = 0.004259
            8'h52: output_q1_11 = 12'h008; // e^(-5.427) = 0.004394
            8'h53: output_q1_11 = 12'h009; // e^(-5.396) = 0.004534
            8'h54: output_q1_11 = 12'h009; // e^(-5.365) = 0.004679
            8'h55: output_q1_11 = 12'h009; // e^(-5.333) = 0.004828
            8'h56: output_q1_11 = 12'h00A; // e^(-5.302) = 0.004982
            8'h57: output_q1_11 = 12'h00A; // e^(-5.271) = 0.005141
            8'h58: output_q1_11 = 12'h00A; // e^(-5.239) = 0.005304
            8'h59: output_q1_11 = 12'h00B; // e^(-5.208) = 0.005473
            8'h5A: output_q1_11 = 12'h00B; // e^(-5.176) = 0.005648
            8'h5B: output_q1_11 = 12'h00B; // e^(-5.145) = 0.005828
            8'h5C: output_q1_11 = 12'h00C; // e^(-5.114) = 0.006014
            8'h5D: output_q1_11 = 12'h00C; // e^(-5.082) = 0.006205
            8'h5E: output_q1_11 = 12'h00D; // e^(-5.051) = 0.006403
            8'h5F: output_q1_11 = 12'h00D; // e^(-5.020) = 0.006607
            8'h60: output_q1_11 = 12'h00D; // e^(-4.988) = 0.006818
            8'h61: output_q1_11 = 12'h00E; // e^(-4.957) = 0.007035
            8'h62: output_q1_11 = 12'h00E; // e^(-4.925) = 0.007259
            8'h63: output_q1_11 = 12'h00F; // e^(-4.894) = 0.007491
            8'h64: output_q1_11 = 12'h00F; // e^(-4.863) = 0.007729
            8'h65: output_q1_11 = 12'h010; // e^(-4.831) = 0.007976
            8'h66: output_q1_11 = 12'h010; // e^(-4.800) = 0.008230
            8'h67: output_q1_11 = 12'h011; // e^(-4.769) = 0.008492
            8'h68: output_q1_11 = 12'h011; // e^(-4.737) = 0.008763
            8'h69: output_q1_11 = 12'h012; // e^(-4.706) = 0.009042
            8'h6A: output_q1_11 = 12'h013; // e^(-4.675) = 0.009330
            8'h6B: output_q1_11 = 12'h013; // e^(-4.643) = 0.009627
            8'h6C: output_q1_11 = 12'h014; // e^(-4.612) = 0.009934
            8'h6D: output_q1_11 = 12'h014; // e^(-4.580) = 0.010251
            8'h6E: output_q1_11 = 12'h015; // e^(-4.549) = 0.010578
            8'h6F: output_q1_11 = 12'h016; // e^(-4.518) = 0.010915
            8'h70: output_q1_11 = 12'h017; // e^(-4.486) = 0.011263
            8'h71: output_q1_11 = 12'h017; // e^(-4.455) = 0.011621
            8'h72: output_q1_11 = 12'h018; // e^(-4.424) = 0.011992
            8'h73: output_q1_11 = 12'h019; // e^(-4.392) = 0.012374
            8'h74: output_q1_11 = 12'h01A; // e^(-4.361) = 0.012768
            8'h75: output_q1_11 = 12'h01A; // e^(-4.329) = 0.013175
            8'h76: output_q1_11 = 12'h01B; // e^(-4.298) = 0.013595
            8'h77: output_q1_11 = 12'h01C; // e^(-4.267) = 0.014028
            8'h78: output_q1_11 = 12'h01D; // e^(-4.235) = 0.014476
            8'h79: output_q1_11 = 12'h01E; // e^(-4.204) = 0.014937
            8'h7A: output_q1_11 = 12'h01F; // e^(-4.173) = 0.015413
            8'h7B: output_q1_11 = 12'h020; // e^(-4.141) = 0.015904
            8'h7C: output_q1_11 = 12'h021; // e^(-4.110) = 0.016411
            8'h7D: output_q1_11 = 12'h022; // e^(-4.078) = 0.016934
            8'h7E: output_q1_11 = 12'h023; // e^(-4.047) = 0.017474
            8'h7F: output_q1_11 = 12'h024; // e^(-4.016) = 0.018031
            8'h80: output_q1_11 = 12'h026; // e^(-3.984) = 0.018605
            8'h81: output_q1_11 = 12'h027; // e^(-3.953) = 0.019198
            8'h82: output_q1_11 = 12'h028; // e^(-3.922) = 0.019810
            8'h83: output_q1_11 = 12'h029; // e^(-3.890) = 0.020441
            8'h84: output_q1_11 = 12'h02B; // e^(-3.859) = 0.021093
            8'h85: output_q1_11 = 12'h02C; // e^(-3.827) = 0.021765
            8'h86: output_q1_11 = 12'h02D; // e^(-3.796) = 0.022459
            8'h87: output_q1_11 = 12'h02F; // e^(-3.765) = 0.023174
            8'h88: output_q1_11 = 12'h030; // e^(-3.733) = 0.023913
            8'h89: output_q1_11 = 12'h032; // e^(-3.702) = 0.024675
            8'h8A: output_q1_11 = 12'h034; // e^(-3.671) = 0.025461
            8'h8B: output_q1_11 = 12'h035; // e^(-3.639) = 0.026273
            8'h8C: output_q1_11 = 12'h037; // e^(-3.608) = 0.027110
            8'h8D: output_q1_11 = 12'h039; // e^(-3.576) = 0.027974
            8'h8E: output_q1_11 = 12'h03B; // e^(-3.545) = 0.028866
            8'h8F: output_q1_11 = 12'h03D; // e^(-3.514) = 0.029786
            8'h90: output_q1_11 = 12'h03E; // e^(-3.482) = 0.030735
            8'h91: output_q1_11 = 12'h040; // e^(-3.451) = 0.031715
            8'h92: output_q1_11 = 12'h043; // e^(-3.420) = 0.032725
            8'h93: output_q1_11 = 12'h045; // e^(-3.388) = 0.033768
            8'h94: output_q1_11 = 12'h047; // e^(-3.357) = 0.034844
            8'h95: output_q1_11 = 12'h049; // e^(-3.325) = 0.035955
            8'h96: output_q1_11 = 12'h04B; // e^(-3.294) = 0.037101
            8'h97: output_q1_11 = 12'h04E; // e^(-3.263) = 0.038283
            8'h98: output_q1_11 = 12'h050; // e^(-3.231) = 0.039503
            8'h99: output_q1_11 = 12'h053; // e^(-3.200) = 0.040762
            8'h9A: output_q1_11 = 12'h056; // e^(-3.169) = 0.042061
            8'h9B: output_q1_11 = 12'h058; // e^(-3.137) = 0.043402
            8'h9C: output_q1_11 = 12'h05B; // e^(-3.106) = 0.044785
            8'h9D: output_q1_11 = 12'h05E; // e^(-3.075) = 0.046212
            8'h9E: output_q1_11 = 12'h061; // e^(-3.043) = 0.047685
            8'h9F: output_q1_11 = 12'h064; // e^(-3.012) = 0.049205
            8'hA0: output_q1_11 = 12'h067; // e^(-2.980) = 0.050773
            8'hA1: output_q1_11 = 12'h06B; // e^(-2.949) = 0.052391
            8'hA2: output_q1_11 = 12'h06E; // e^(-2.918) = 0.054061
            8'hA3: output_q1_11 = 12'h072; // e^(-2.886) = 0.055784
            8'hA4: output_q1_11 = 12'h075; // e^(-2.855) = 0.057561
            8'hA5: output_q1_11 = 12'h079; // e^(-2.824) = 0.059396
            8'hA6: output_q1_11 = 12'h07D; // e^(-2.792) = 0.061289
            8'hA7: output_q1_11 = 12'h081; // e^(-2.761) = 0.063242
            8'hA8: output_q1_11 = 12'h085; // e^(-2.729) = 0.065258
            8'hA9: output_q1_11 = 12'h089; // e^(-2.698) = 0.067337
            8'hAA: output_q1_11 = 12'h08E; // e^(-2.667) = 0.069483
            8'hAB: output_q1_11 = 12'h092; // e^(-2.635) = 0.071698
            8'hAC: output_q1_11 = 12'h097; // e^(-2.604) = 0.073983
            8'hAD: output_q1_11 = 12'h09C; // e^(-2.573) = 0.076341
            8'hAE: output_q1_11 = 12'h0A1; // e^(-2.541) = 0.078774
            8'hAF: output_q1_11 = 12'h0A6; // e^(-2.510) = 0.081284
            8'hB0: output_q1_11 = 12'h0AB; // e^(-2.478) = 0.083875
            8'hB1: output_q1_11 = 12'h0B1; // e^(-2.447) = 0.086548
            8'hB2: output_q1_11 = 12'h0B6; // e^(-2.416) = 0.089306
            8'hB3: output_q1_11 = 12'h0BC; // e^(-2.384) = 0.092152
            8'hB4: output_q1_11 = 12'h0C2; // e^(-2.353) = 0.095089
            8'hB5: output_q1_11 = 12'h0C8; // e^(-2.322) = 0.098120
            8'hB6: output_q1_11 = 12'h0CF; // e^(-2.290) = 0.101247
            8'hB7: output_q1_11 = 12'h0D5; // e^(-2.259) = 0.104473
            8'hB8: output_q1_11 = 12'h0DC; // e^(-2.227) = 0.107803
            8'hB9: output_q1_11 = 12'h0E3; // e^(-2.196) = 0.111239
            8'hBA: output_q1_11 = 12'h0EB; // e^(-2.165) = 0.114784
            8'hBB: output_q1_11 = 12'h0F2; // e^(-2.133) = 0.118442
            8'hBC: output_q1_11 = 12'h0FA; // e^(-2.102) = 0.122217
            8'hBD: output_q1_11 = 12'h102; // e^(-2.071) = 0.126112
            8'hBE: output_q1_11 = 12'h10A; // e^(-2.039) = 0.130131
            8'hBF: output_q1_11 = 12'h113; // e^(-2.008) = 0.134278
            8'hC0: output_q1_11 = 12'h11B; // e^(-1.976) = 0.138557
            8'hC1: output_q1_11 = 12'h124; // e^(-1.945) = 0.142973
            8'hC2: output_q1_11 = 12'h12E; // e^(-1.914) = 0.147530
            8'hC3: output_q1_11 = 12'h137; // e^(-1.882) = 0.152231
            8'hC4: output_q1_11 = 12'h141; // e^(-1.851) = 0.157083
            8'hC5: output_q1_11 = 12'h14B; // e^(-1.820) = 0.162089
            8'hC6: output_q1_11 = 12'h156; // e^(-1.788) = 0.167255
            8'hC7: output_q1_11 = 12'h161; // e^(-1.757) = 0.172585
            8'hC8: output_q1_11 = 12'h16C; // e^(-1.725) = 0.178086
            8'hC9: output_q1_11 = 12'h178; // e^(-1.694) = 0.183761
            8'hCA: output_q1_11 = 12'h184; // e^(-1.663) = 0.189618
            8'hCB: output_q1_11 = 12'h190; // e^(-1.631) = 0.195661
            8'hCC: output_q1_11 = 12'h19D; // e^(-1.600) = 0.201897
            8'hCD: output_q1_11 = 12'h1AA; // e^(-1.569) = 0.208331
            8'hCE: output_q1_11 = 12'h1B8; // e^(-1.537) = 0.214970
            8'hCF: output_q1_11 = 12'h1C6; // e^(-1.506) = 0.221821
            8'hD0: output_q1_11 = 12'h1D4; // e^(-1.475) = 0.228891
            8'hD1: output_q1_11 = 12'h1E3; // e^(-1.443) = 0.236186
            8'hD2: output_q1_11 = 12'h1F3; // e^(-1.412) = 0.243713
            8'hD3: output_q1_11 = 12'h203; // e^(-1.380) = 0.251480
            8'hD4: output_q1_11 = 12'h213; // e^(-1.349) = 0.259495
            8'hD5: output_q1_11 = 12'h224; // e^(-1.318) = 0.267765
            8'hD6: output_q1_11 = 12'h235; // e^(-1.286) = 0.276298
            8'hD7: output_q1_11 = 12'h247; // e^(-1.255) = 0.285104
            8'hD8: output_q1_11 = 12'h25A; // e^(-1.224) = 0.294190
            8'hD9: output_q1_11 = 12'h26D; // e^(-1.192) = 0.303566
            8'hDA: output_q1_11 = 12'h281; // e^(-1.161) = 0.313240
            8'hDB: output_q1_11 = 12'h295; // e^(-1.129) = 0.323223
            8'hDC: output_q1_11 = 12'h2AB; // e^(-1.098) = 0.333524
            8'hDD: output_q1_11 = 12'h2C0; // e^(-1.067) = 0.344154
            8'hDE: output_q1_11 = 12'h2D7; // e^(-1.035) = 0.355122
            8'hDF: output_q1_11 = 12'h2EE; // e^(-1.004) = 0.366440
            8'hE0: output_q1_11 = 12'h306; // e^(-0.973) = 0.378118
            8'hE1: output_q1_11 = 12'h31F; // e^(-0.941) = 0.390169
            8'hE2: output_q1_11 = 12'h338; // e^(-0.910) = 0.402603
            8'hE3: output_q1_11 = 12'h352; // e^(-0.878) = 0.415434
            8'hE4: output_q1_11 = 12'h36D; // e^(-0.847) = 0.428674
            8'hE5: output_q1_11 = 12'h389; // e^(-0.816) = 0.442336
            8'hE6: output_q1_11 = 12'h3A6; // e^(-0.784) = 0.456433
            8'hE7: output_q1_11 = 12'h3C4; // e^(-0.753) = 0.470979
            8'hE8: output_q1_11 = 12'h3E3; // e^(-0.722) = 0.485989
            8'hE9: output_q1_11 = 12'h403; // e^(-0.690) = 0.501478
            8'hEA: output_q1_11 = 12'h423; // e^(-0.659) = 0.517460
            8'hEB: output_q1_11 = 12'h445; // e^(-0.627) = 0.533951
            8'hEC: output_q1_11 = 12'h468; // e^(-0.596) = 0.550968
            8'hED: output_q1_11 = 12'h48C; // e^(-0.565) = 0.568527
            8'hEE: output_q1_11 = 12'h4B1; // e^(-0.533) = 0.586646
            8'hEF: output_q1_11 = 12'h4D7; // e^(-0.502) = 0.605343
            8'hF0: output_q1_11 = 12'h4FF; // e^(-0.471) = 0.624635
            8'hF1: output_q1_11 = 12'h528; // e^(-0.439) = 0.644542
            8'hF2: output_q1_11 = 12'h552; // e^(-0.408) = 0.665083
            8'hF3: output_q1_11 = 12'h57D; // e^(-0.376) = 0.686279
            8'hF4: output_q1_11 = 12'h5AA; // e^(-0.345) = 0.708151
            8'hF5: output_q1_11 = 12'h5D8; // e^(-0.314) = 0.730720
            8'hF6: output_q1_11 = 12'h608; // e^(-0.282) = 0.754008
            8'hF7: output_q1_11 = 12'h639; // e^(-0.251) = 0.778038
            8'hF8: output_q1_11 = 12'h66C; // e^(-0.220) = 0.802834
            8'hF9: output_q1_11 = 12'h6A0; // e^(-0.188) = 0.828420
            8'hFA: output_q1_11 = 12'h6D6; // e^(-0.157) = 0.854821
            8'hFB: output_q1_11 = 12'h70E; // e^(-0.125) = 0.882064
            8'hFC: output_q1_11 = 12'h748; // e^(-0.094) = 0.910176
            8'hFD: output_q1_11 = 12'h783; // e^(-0.063) = 0.939183
            8'hFE: output_q1_11 = 12'h7C0; // e^(-0.031) = 0.969114
            8'hFF: output_q1_11 = 12'h800; // e^(0.000) = 1.000000
            default: output_q1_11 = 12'h000;
        endcase
    end

endmodule
